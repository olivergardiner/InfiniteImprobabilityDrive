Inifinite Improbability Drive

VIN 21  0    DC 0    AC 1 SIN(0 0.7 1K)
VDD 50  0    DC 10   AC 0
VB  40  0    DC 5    AC 0
VDX 51  0    DC 10   AC 0
VDY 52  0    DC 10   AC 0

.INCLUDE OPAMP1.cir

.MODEL J201 NJF(Beta=1.621m Betatce=-500m Rd=1 Rs=1 Lambda=2.236m Vto=-600m Vtotc=-2.5m Is=114.5f Cgd=4.667p M=227.1m Pb=500m Fc=500m Cgs=2.992p Kf=0.6042f Af=1)
.MODEL J202 NJF(Beta=985.5u Betatce=-500m Rd=1 Rs=1 Lambda=7m Vto=-1.612 Vtotc=-2.5m Is=114.5f Xti=3 Cgd=4.667p M=227.1m Pb=500m Fc=500m Cgs=2.992p Kf=0.3604f Af=1)
.MODEL 2N5088 NPN(IS=5.911f ISE=5.911f ISC=0 XTI=3 BF=1122 BR=1.271 IKF=14.92m IKR=0 XTB=1.5 VAF=62.37 VAR=21.5 VJE=0.65 VJC=0.65 RE=0.15 RC=1.61 RB=10 CJE=4.973p CJC=4.017p XCJC=0.75 FC=0.5 NF=1 NR=1 NE=1.394 NC=2 MJE=0.4146 MJC=0.3174 TF=821.7p TR=4.673n ITF=0.35 VTF=4 XTF=7 EG=1.11 VCEO=35 ICRATING=50m MFG=NSC)
.MODEL 2N5086 PNP(IS=28.000f ISE=24.903f ISC=0.125p XTI=3.300 BF=284.436 BR=4.800 IKF=0.380 IKR=0.932 XTB=1.600 VAF=43.0 VAR=6.960 VJE=1.0 VJC=0.900 RE=0.300 RC=2.251 RB=2.200 RBM=1.500 IRB=0.100m CJE=11.800p CJC=8.700p XCJC=0.650 FC=0.750 NF=1.0 NR=1.005 NE=2.234 NC=2.074 MJE=0.435 MJC=0.600 TF=0.600n TR=2.604n PTF=1.0 ITF=0.314 VTF=2.0 XTF=6.500 EG=1.110 VCEO=50 ICRATING=50m MFG=SIEMENS)
.MODEL 1N4148 D(Is=2.52n Rs=.568 N=1.752 Cjo=4p M=.4 tt=20n)

C8  21 22    47N
J6  24 22 23 J201
R14 22 40    470K
R15  0 22    270K
R8   0 23    51K
R10 24 50    47K
C9  24 25    47N
R17  0 25    680K
R9   0 26    6.8K
C13  0 28    47N
R18  0 32    680K
C12 23 32    4.7N
J8  27 25 26 J201
J9  28 32 26 J201
Q2  27 27 51 2N5086
Q3  28 28 52 2N5086

Q4  29 27 50 2N5086
Q6  29 29  0 2N5088
Q5  31 28 50 2N5086
Q7  30 29  0 2N5088
R16 30 40    4.7K
R32 31 40    4.7K

RV  25 32    1000K

R19 30 34    220K
R21 31 34    220K
R20 34 35    220K
X1  40 34 35 OPAMP1

RL   0 35    100K

*.OPTIONS NOACCT RELTOL=.01
.OPTIONS NOACCT
.TRAN 10US 50MS 45MS

.END